library ieee;
use ieee.std_logic_1164.all;

entity part1 is
	port(address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		clock : IN STD_LOGIC := '1';
		data : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		wren : IN STD_LOGIC ;
		q : OUT STD_LOGIC_VECTOR (3 DOWNTO 0) );
end part1;

architecture be of part1 is
	
	component ram32x4
		PORT ( address : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
				clock : IN STD_LOGIC := '1';
				data : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
				wren : IN STD_LOGIC ;
				q : OUT STD_LOGIC_VECTOR (3 DOWNTO 0) );
	end component;
	
begin

	inst1: ram32x4
	port map(address => address,
				clock => clock,
				data => data,
				wren => wren,
				q => q);

end be;